LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
 
LIBRARY WORK;
USE WORK.HdmiPkg.ALL;

PACKAGE GamePkg IS
  CONSTANT c_GAME_SCALE : INTEGER := 20;
  
  CONSTANT c_REFRESH_RATE : INTEGER := c_PIXEL_CLK_FREQ/c_GAME_SCALE;
  CONSTANT c_GAME_WIDTH : INTEGER := c_FRAME_WIDTH/c_GAME_SCALE;
  CONSTANT c_GAME_HEIGHT : INTEGER := c_FRAME_HEIGHT/c_GAME_SCALE;
 
  -- CONSTANT c_SCORE_LIMIT : INTEGER := 100;
  -- CONSTANT c_SCORE_WIDTH : INTEGER := 3;
  -- CONSTANT c_SCORE_HEIGHT : INTEGER := 5;
  -- CONSTANT c_SCORE_Y_POS : INTEGER := 1;
  -- CONSTANT c_SCORE_COL : INTEGER := c_GAME_WIDTH - 3*c_SCORE_WIDTH;
   
  CONSTANT c_MIN_SNAKE_SIZE : INTEGER := 3;
  CONSTANT c_MAX_SNAKE_SIZE : INTEGER := 10;
  
  CONSTANT c_SNAKE_SPEED : INTEGER := c_REFRESH_RATE; 
END PACKAGE GamePkg; 