LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

PACKAGE HdmiPkg IS 
    CONSTANT c_HDMI_CLK_FREQ : INTEGER := 400000000;
    CONSTANT c_PIXEL_CLK_FREQ : INTEGER := c_HDMI_CLK_FREQ/10;

    SUBTYPE t_Byte IS STD_LOGIC_VECTOR(7 DOWNTO 0);
    SUBTYPE t_RGB IS STD_LOGIC_VECTOR(23 DOWNTO 0); 
    
    -- Timing parameters for 800x600@60Hz
    CONSTANT c_FRAME_WIDTH_800x600   : INTEGER := 800;
    CONSTANT c_H_FRONT_PORCH_800x600 : INTEGER := 40;
    CONSTANT c_H_BACK_PORCH_800x600  : INTEGER := 88;
    CONSTANT c_H_PULSE_WIDTH_800x600 : INTEGER := 128;
    CONSTANT c_FRAME_HEIGHT_800x600  : INTEGER := 600;
    CONSTANT c_V_FRONT_PORCH_800x600 : INTEGER := 1;
    CONSTANT c_V_BACK_PORCH_800x600  : INTEGER := 23;
    CONSTANT c_V_PULSE_WIDTH_800x600 : INTEGER := 4;
    
    -- Timing parameters for 640x480@60Hz
    CONSTANT c_FRAME_WIDTH_640x480   : INTEGER := 640;
    CONSTANT c_H_FRONT_PORCH_640x480 : INTEGER := 16;
    CONSTANT c_H_BACK_PORCH_640x480  : INTEGER := 48;
    CONSTANT c_H_PULSE_WIDTH_640x480 : INTEGER := 96;
    CONSTANT c_FRAME_HEIGHT_640x480  : INTEGER := 480;
    CONSTANT c_V_FRONT_PORCH_640x480 : INTEGER := 10;
    CONSTANT c_V_BACK_PORCH_640x480  : INTEGER := 33;
    CONSTANT c_V_PULSE_WIDTH_640x480 : INTEGER := 2;
    
    CONSTANT c_FRAME_WIDTH   : INTEGER := c_FRAME_WIDTH_800x600;
    CONSTANT c_H_FRONT_PORCH : INTEGER := c_H_FRONT_PORCH_800x600;
    CONSTANT c_H_BACK_PORCH  : INTEGER := c_H_BACK_PORCH_800x600;
    CONSTANT c_H_PULSE_WIDTH : INTEGER := c_H_PULSE_WIDTH_800x600;
    CONSTANT c_H_BLANK       : INTEGER := c_H_FRONT_PORCH + c_H_BACK_PORCH + c_H_PULSE_WIDTH;
    
    CONSTANT c_FRAME_HEIGHT  : INTEGER := c_FRAME_HEIGHT_800x600;
    CONSTANT c_V_FRONT_PORCH : INTEGER := c_V_FRONT_PORCH_800x600;
    CONSTANT c_V_BACK_PORCH  : INTEGER := c_V_BACK_PORCH_800x600;
    CONSTANT c_V_PULSE_WIDTH : INTEGER := c_V_PULSE_WIDTH_800x600;
    CONSTANT c_V_BLANK       : INTEGER := c_V_FRONT_PORCH + c_V_BACK_PORCH + c_V_PULSE_WIDTH;
    
    CONSTANT c_H_MAX : INTEGER := c_FRAME_WIDTH + c_H_BLANK;
    CONSTANT c_V_MAX : INTEGER := c_FRAME_HEIGHT + c_V_BLANK;
	
	CONSTANT c_DISPLAY_RESOLUTION : INTEGER := c_FRAME_WIDTH * c_FRAME_HEIGHT;
	CONSTANT c_MAX_RESOLUTION : INTEGER := c_H_MAX * c_V_MAX; 
END HdmiPkg;
