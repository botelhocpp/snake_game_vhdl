LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
 
LIBRARY WORK;
USE WORK.HdmiPkg.ALL;

PACKAGE GamePkg IS
  CONSTANT c_GAME_SCALE : INTEGER := 20;
  CONSTANT c_REFRESH_RATE : INTEGER := c_PIXEL_CLK_FREQ/c_GAME_SCALE;

  CONSTANT c_GAME_WIDTH : INTEGER := c_FRAME_WIDTH/c_GAME_SCALE;
  CONSTANT c_GAME_HEIGHT : INTEGER := c_FRAME_HEIGHT/c_GAME_SCALE;

  CONSTANT c_GAME_X_MIDDLE  : INTEGER := c_GAME_WIDTH/2 - 1;
  CONSTANT c_GAME_Y_MIDDLE  : INTEGER := c_GAME_HEIGHT/2 - 1;

  -- Game limits
  CONSTANT c_GAME_LIMIT_LEFT_LINE : INTEGER := 1;
  CONSTANT c_GAME_LIMIT_RIGHT_LINE : INTEGER := c_GAME_WIDTH - 2;
  CONSTANT c_GAME_LIMIT_UPPER_LINE : INTEGER := 1;
  CONSTANT c_GAME_LIMIT_LOWER_LINE : INTEGER := c_GAME_HEIGHT - 2;

  -- Game valid positions
  CONSTANT c_GAME_FIRST_COL : INTEGER := c_GAME_LIMIT_LEFT_LINE + 1;
  CONSTANT c_GAME_LAST_COL : INTEGER := c_GAME_LIMIT_RIGHT_LINE - 1;
  CONSTANT c_GAME_FIRST_ROW : INTEGER := c_GAME_LIMIT_UPPER_LINE + 1;
  CONSTANT c_GAME_LAST_ROW : INTEGER := c_GAME_LIMIT_LOWER_LINE - 1;
 
  -- Snake dimensions and position
  -- CONSTANT c_SCORE_LIMIT : INTEGER := 999;
  -- CONSTANT c_SCORE_WIDTH : INTEGER := 3;
  -- CONSTANT c_SCORE_HEIGHT : INTEGER := 5;
  -- CONSTANT c_SCORE_Y_POS : INTEGER := c_GAME_LIMIT_UPPER_LINE + 2;
  -- CONSTANT c_SCORE_COL : INTEGER := c_GAME_WIDTH - 3*c_SCORE_WIDTH;
   
  CONSTANT c_MIN_SNAKE_SIZE : INTEGER := 3;
  CONSTANT c_MAX_SNAKE_SIZE : INTEGER := 10; -- c_GAME_WIDTH * c_GAME_HEIGHT;
  
  CONSTANT c_MAX_SNAKE_SPEED : INTEGER := 2*c_REFRESH_RATE; 
  CONSTANT c_SNAKE_SPEED_EASY : INTEGER := 2*c_REFRESH_RATE; 
  CONSTANT c_SNAKE_SPEED_NORMAL : INTEGER := c_REFRESH_RATE; 
  CONSTANT c_SNAKE_SPEED_HARD : INTEGER := c_REFRESH_RATE/2; 
END PACKAGE GamePkg; 